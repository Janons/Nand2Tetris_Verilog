module and( 
    input a, 
    input b, 
    output out );

    assing out = a&b;
endmodule