# ifndef or_n2t