


module not (in , out);
    input in;
    output out;

    //module code goes here
    nand result(in , in , out);

    
endmodule