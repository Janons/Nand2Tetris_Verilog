# ifndef or_n2t


module not (a,b, in);

    wire nand_a_b

    nand nand_b_a(nand_a_b, a ,b)
    not_n2t and_n2t(nand_a_b,out)

    //module code goes here
    nand result(a , b , out);

    
endmodule