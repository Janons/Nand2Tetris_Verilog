module top_module ( input a, input b, output out );
    mod_a inst(a,b,out);
endmodule